`timescale 1ns / 1ps

module control_unit();
endmodule
